module execute();

`include "funcs.v"

endmodule
