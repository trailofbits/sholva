module alu(
  input [8:0] cntl,
  input [31:0] opnd0_r,
  input [31:0] opnd1_r
);

// TODO: extend operands to 33 bits for carries, mix in carry bit from EFLAGS when
// requested

endmodule
