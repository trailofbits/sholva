module circuit(
input [1237:0] current,
input [1237:0] next,

output [0:0] result
);
wire In_error_flag = current[0: 0];
wire In_register_AF = current[121: 121];
wire In_register_CF = current[122: 122];
wire [31:0] In_register_CSBASE = current[154: 123];
wire [7:0] In_register_DF = current[162: 155];
wire [31:0] In_register_DSBASE = current[194: 163];
wire [31:0] In_register_EAX = current[226: 195];
wire [31:0] In_register_EBP = current[258: 227];
wire [31:0] In_register_EBX = current[290: 259];
wire [31:0] In_register_ECX = current[322: 291];
wire [31:0] In_register_EDI = current[354: 323];
wire [31:0] In_register_EDX = current[386: 355];
wire [31:0] In_register_EIP = current[418: 387];
wire [31:0] In_register_ESBASE = current[450: 419];
wire [31:0] In_register_ESI = current[482: 451];
wire [31:0] In_register_ESP = current[514: 483];
wire [31:0] In_register_FSBASE = current[546: 515];
wire [31:0] In_register_GSBASE = current[578: 547];
wire In_register_OF = current[579: 579];
wire In_register_PF = current[580: 580];
wire In_register_SF = current[581: 581];
wire [31:0] In_register_SSBASE = current[613: 582];
wire In_register_ZF = current[614: 614];
wire [63:0] In_timestamp = current[678: 615];
wire Out_error_flag = next[0: 0];
wire Out_register_AF = next[121: 121];
wire Out_register_CF = next[122: 122];
wire [31:0] Out_register_CSBASE = next[154: 123];
wire [7:0] Out_register_DF = next[162: 155];
wire [31:0] Out_register_DSBASE = next[194: 163];
wire [31:0] Out_register_EAX = next[226: 195];
wire [31:0] Out_register_EBP = next[258: 227];
wire [31:0] Out_register_EBX = next[290: 259];
wire [31:0] Out_register_ECX = next[322: 291];
wire [31:0] Out_register_EDI = next[354: 323];
wire [31:0] Out_register_EDX = next[386: 355];
wire [31:0] Out_register_EIP = next[418: 387];
wire [31:0] Out_register_ESBASE = next[450: 419];
wire [31:0] Out_register_ESI = next[482: 451];
wire [31:0] Out_register_ESP = next[514: 483];
wire [31:0] Out_register_FSBASE = next[546: 515];
wire [31:0] Out_register_GSBASE = next[578: 547];
wire Out_register_OF = next[579: 579];
wire Out_register_PF = next[580: 580];
wire Out_register_SF = next[581: 581];
wire [31:0] Out_register_SSBASE = next[613: 582];
wire Out_register_ZF = next[614: 614];
wire [63:0] Out_timestamp = next[678: 615];
wire [119:0] instruction_bits = current[120: 1];
wire [7:0] vf = 8'b00010001;
wire [7:0] v114 = instruction_bits[7: 0];
wire v115 = vf == v114;
wire [1:0] v10 = 2'b11;
wire [1:0] v116 = instruction_bits[15: 14];
wire v117 = v10 == v116;
wire [103:0] v11 = 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
wire [103:0] v118 = instruction_bits[119: 16];
wire v119 = v11 == v118;
wire v11a = v115 & v117 & v119;
wire v11b = v11a;
wire v11c = v11b;
wire [2:0] v125 = instruction_bits[10: 8];
wire [2:0] v16c = { v125 };
wire [2:0] v6 = 3'b000;
wire v16d = v16c == v6;
wire v16e = v16d;
wire v16f = v11a & v16e;
wire v185 = v16f;
wire [2:0] v13d = instruction_bits[13: 11];
wire [2:0] v13e = { v13d };
wire v13a = 1'b1;
wire [2:0] v139 = ( v11c ) ? v13e : v6;
wire [31:0] v13c = ( v139 == 3'd0) ? In_register_EAX : 
	( v139 == 3'd1) ? In_register_ECX : 
	( v139 == 3'd2) ? In_register_EDX : 
	( v139 == 3'd3) ? In_register_EBX : 
	( v139 == 3'd4) ? In_register_ESP : 
	( v139 == 3'd5) ? In_register_EBP : 
	( v139 == 3'd6) ? In_register_ESI : In_register_EDI;
wire [31:0] v150 = v13c;
wire [2:0] v126 = { v125 };
wire v122 = 1'b1;
wire [2:0] v121 = ( v11c ) ? v126 : v6;
wire [31:0] v124 = ( v121 == 3'd0) ? In_register_EAX : 
	( v121 == 3'd1) ? In_register_ECX : 
	( v121 == 3'd2) ? In_register_EDX : 
	( v121 == 3'd3) ? In_register_EBX : 
	( v121 == 3'd4) ? In_register_ESP : 
	( v121 == 3'd5) ? In_register_EBP : 
	( v121 == 3'd6) ? In_register_ESI : In_register_EDI;
wire [31:0] v138 = v124;
wire [31:0] v152 = v150 + v138;
wire [7:0] v11d = { 7'b0000000, In_register_CF };
wire [31:0] v151 = { 24'b000000000000000000000000, v11d };
wire [31:0] v153 = v152 + v151;
wire ve = 1'b1;
wire [31:0] v188 = ( v185 ) ? v153 : In_register_EAX;
wire [31:0] v1a9 = v188;
wire v1aa = v1a9 == Out_register_EAX;
wire [2:0] v8 = 3'b011;
wire v173 = v16c == v8;
wire v174 = v173;
wire v175 = v11a & v174;
wire v189 = v175;
wire [31:0] v18c = ( v189 ) ? v153 : In_register_EBX;
wire [31:0] v1ac = v18c;
wire v1ad = v1ac == Out_register_EBX;
wire [2:0] va = 3'b111;
wire v179 = v16c == va;
wire v17a = v179;
wire v17b = v11a & v17a;
wire v199 = v17b;
wire [31:0] v19c = ( v199 ) ? v153 : In_register_EDI;
wire [31:0] v1b8 = v19c;
wire v1b9 = v1b8 == Out_register_EDI;
wire [7:0] v15c = v153[7:0];
wire [2:0] v15d_aux = v15c[0] + v15c[1] + v15c[2] + v15c[3] + v15c[4] + v15c[5] + v15c[6] + v15c[7];
wire v15d = { 5'b00000, v15d_aux };
wire [7:0] v13 = 8'b00000001;
wire [7:0] v15e = v15d & v13;
wire [7:0] v15f = v15e ^ v13;
wire v1a7 = v15f[0:0];
wire v1e3 = v1a7;
wire v1e4 = v1e3 == Out_register_PF;
wire [2:0] vb = 3'b010;
wire v17c = v16c == vb;
wire v17d = v17c;
wire v17e = v11a & v17d;
wire v191 = v17e;
wire [31:0] v194 = ( v191 ) ? v153 : In_register_EDX;
wire [31:0] v1b2 = v194;
wire v1b3 = v1b2 == Out_register_EDX;
wire [2:0] vc = 3'b110;
wire v17f = v16c == vc;
wire v180 = v17f;
wire v181 = v11a & v180;
wire v195 = v181;
wire [31:0] v198 = ( v195 ) ? v153 : In_register_ESI;
wire [31:0] v1b5 = v198;
wire v1b6 = v1b5 == Out_register_ESI;
wire [63:0] v2 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
wire [63:0] v1c = In_timestamp + v2;
wire v1d = v1c == Out_timestamp;
wire [31:0] v1d0 = In_register_GSBASE;
wire v1d1 = v1d0 == Out_register_GSBASE;
wire [31:0] v15 = 32'b00000000000000000000000000000000;
wire v165 = v153 == v15;
wire v1e9 = v165;
wire v1ea = v1e9 == Out_register_ZF;
wire [31:0] v1c7 = In_register_SSBASE;
wire v1c8 = v1c7 == Out_register_SSBASE;
wire [2:0] vd = 3'b100;
wire v182 = v16c == vd;
wire v183 = v182;
wire v184 = v11a & v183;
wire v19d = v184;
wire [31:0] v1a0 = ( v19d ) ? v153 : In_register_ESP;
wire [31:0] v1bb = v1a0;
wire v1bc = v1bb == Out_register_ESP;
wire [31:0] v12 = 32'b00000000000000000000000000000010;
wire [31:0] v11f = v12;
wire [31:0] v120 = In_register_EIP + v11f;
wire [31:0] v1c1 = v120;
wire v1c2 = v1c1 == Out_register_EIP;
wire [2:0] v7 = 3'b101;
wire v170 = v16c == v7;
wire v171 = v170;
wire v172 = v11a & v171;
wire v1a1 = v172;
wire [31:0] v1a4 = ( v1a1 ) ? v153 : In_register_EBP;
wire [31:0] v1be = v1a4;
wire v1bf = v1be == Out_register_EBP;
wire [31:0] v1c4 = In_register_CSBASE;
wire v1c5 = v1c4 == Out_register_CSBASE;
wire [31:0] v1ca = In_register_ESBASE;
wire v1cb = v1ca == Out_register_ESBASE;
wire [31:0] v1cd = In_register_DSBASE;
wire v1ce = v1cd == Out_register_DSBASE;
wire [2:0] v9 = 3'b001;
wire v176 = v16c == v9;
wire v177 = v176;
wire v178 = v11a & v177;
wire v18d = v178;
wire [31:0] v190 = ( v18d ) ? v153 : In_register_ECX;
wire [31:0] v1af = v190;
wire v1b0 = v1af == Out_register_ECX;
wire [31:0] v1d3 = In_register_FSBASE;
wire v1d4 = v1d3 == Out_register_FSBASE;
wire [31:0] v160 = v153 ^ v150;
wire [31:0] v161 = v160 ^ v138;
wire [7:0] v162 = v161[7:0];
wire [7:0] v14 = 8'b00000100;
wire [7:0] v163 = v162 >> v14;
wire [7:0] v164 = v163 & v13;
wire v1a5 = v164[0:0];
wire v1d6 = v1a5;
wire v1d7 = v1d6 == Out_register_AF;
wire v166 = $signed(v153) < $signed(v15);
wire v1e6 = v166;
wire v1e7 = v1e6 == Out_register_SF;
wire v1eb = In_error_flag == Out_error_flag;
wire v154 = v152 < v138;
wire v155 = v152 < v150;
wire v156 = v154 | v155;
wire v157 = v153 < v152;
wire v158 = v153 < v151;
wire v159 = v157 | v158;
wire [7:0] v15a = { 7'b0000000, v159 };
wire [7:0] v15b = ( v156 == 1'd0) ? v15a : v13;
wire v1a6 = v15b[0:0];
wire v1d9 = v1a6;
wire v1da = v1d9 == Out_register_CF;
wire [7:0] v1dc = In_register_DF;
wire v1dd = v1dc == Out_register_DF;
wire v1de = v1dd;
wire [31:0] v167 = v153 ^ v138;
wire [31:0] v16 = 32'b00000000000000000000000000011111;
wire [31:0] v168 = v167 >> v16;
wire [31:0] v169 = v160 >> v16;
wire [31:0] v16a = v168 + v169;
wire v16b = v16a == v12;
wire v1e0 = v16b;
wire v1e1 = v1e0 == Out_register_OF;
wire v1ec = v1aa & v1ad & v1b9 & v1e4 & v1b3 & v1b6 & v11c & v1d & v1d1 & v1ea & v1c8 & v1bc & v1c2 & v1bf & v1c5 & v1cb & v1ce & v1b0 & v1d4 & v1d7 & v1e7 & v1eb & v1da & v1de & v1e1;
wire [7:0] v17 = 8'b11111001;
wire v1ed = v17 == v114;
wire [111:0] v18 = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
wire [111:0] v1ee = instruction_bits[119: 8];
wire v1ef = v18 == v1ee;
wire v1f0 = v1ed & v1ef;
wire v1f1 = v1f0;
wire v1f2 = v1f1;
wire [31:0] v1fa = In_register_EBX;
wire v1fb = v1fa == Out_register_EBX;
wire [31:0] v206 = In_register_EDI;
wire v207 = v206 == Out_register_EDI;
wire [31:0] v221 = In_register_FSBASE;
wire v222 = v221 == Out_register_FSBASE;
wire v231 = In_register_PF;
wire v232 = v231 == Out_register_PF;
wire [31:0] v203 = In_register_ESI;
wire v204 = v203 == Out_register_ESI;
wire v239 = In_error_flag == Out_error_flag;
wire [31:0] v20c = In_register_EBP;
wire v20d = v20c == Out_register_EBP;
wire v22e = In_register_OF;
wire v22f = v22e == Out_register_OF;
wire [31:0] v212 = In_register_CSBASE;
wire v213 = v212 == Out_register_CSBASE;
wire [31:0] v1fd = In_register_ECX;
wire v1fe = v1fd == Out_register_ECX;
wire [31:0] v209 = In_register_ESP;
wire v20a = v209 == Out_register_ESP;
wire v227 = ve;
wire v228 = v227 == Out_register_CF;
wire [7:0] v22a = In_register_DF;
wire v22b = v22a == Out_register_DF;
wire v22c = v22b;
wire v234 = In_register_SF;
wire v235 = v234 == Out_register_SF;
wire [31:0] v215 = In_register_SSBASE;
wire v216 = v215 == Out_register_SSBASE;
wire [31:0] v19 = 32'b00000000000000000000000000000001;
wire [31:0] v1f4 = v19;
wire [31:0] v1f5 = In_register_EIP + v1f4;
wire [31:0] v20f = v1f5;
wire v210 = v20f == Out_register_EIP;
wire [31:0] v218 = In_register_ESBASE;
wire v219 = v218 == Out_register_ESBASE;
wire [31:0] v21b = In_register_DSBASE;
wire v21c = v21b == Out_register_DSBASE;
wire [31:0] v200 = In_register_EDX;
wire v201 = v200 == Out_register_EDX;
wire [31:0] v21e = In_register_GSBASE;
wire v21f = v21e == Out_register_GSBASE;
wire v224 = In_register_AF;
wire v225 = v224 == Out_register_AF;
wire [31:0] v1f7 = In_register_EAX;
wire v1f8 = v1f7 == Out_register_EAX;
wire v237 = In_register_ZF;
wire v238 = v237 == Out_register_ZF;
wire v23a = v1fb & v207 & v1d & v1f2 & v222 & v232 & v204 & v239 & v20d & v22f & v213 & v1fe & v20a & v228 & v22c & v235 & v216 & v210 & v219 & v21c & v201 & v21f & v225 & v1f8 & v238;
wire [4:0] v3 = 5'b10111;
wire [4:0] v1e = instruction_bits[7: 3];
wire v1f = v3 == v1e;
wire [79:0] v4 = 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
wire [79:0] v20 = instruction_bits[119: 40];
wire v21 = v4 == v20;
wire v22 = v1f & v21;
wire v23 = v3 == v1e;
wire v24 = v4 == v20;
wire v25 = v23 & v24;
wire v26 = v3 == v1e;
wire v27 = v4 == v20;
wire v28 = v26 & v27;
wire v29 = v22 | v25 | v28;
wire v2a = v29;
wire v101 = In_register_OF;
wire v103 = v101 == Out_register_OF;
wire [2:0] v4b = instruction_bits[2: 0];
wire [2:0] v4c = { v4b };
wire v53 = v4c == v8;
wire v54 = v53;
wire v55 = v22 & v54;
wire [2:0] v65 = { v4b };
wire v6c = v65 == v8;
wire v6d = v6c;
wire v6e = v25 & v6d;
wire [2:0] v7e = { v4b };
wire v85 = v7e == v8;
wire v86 = v85;
wire v87 = v28 & v86;
wire v9b = v55 | v6e | v87;
wire [31:0] v46 = instruction_bits[39: 8];
wire [31:0] v4a = ( v22 | v25 ) ? v46 : v46;
wire [31:0] v9e = ( v9b ) ? v4a : In_register_EBX;
wire [31:0] vbc = v9e;
wire vbe = vbc == Out_register_EBX;
wire v109 = In_register_SF;
wire v10b = v109 == Out_register_SF;
wire v56 = v4c == v9;
wire v57 = v56;
wire v58 = v22 & v57;
wire v6f = v65 == v9;
wire v70 = v6f;
wire v71 = v25 & v70;
wire v88 = v7e == v9;
wire v89 = v88;
wire v8a = v28 & v89;
wire v9f = v58 | v71 | v8a;
wire [31:0] va2 = ( v9f ) ? v4a : In_register_ECX;
wire [31:0] vc0 = va2;
wire vc2 = vc0 == Out_register_ECX;
wire v5f = v4c == vc;
wire v60 = v5f;
wire v61 = v22 & v60;
wire v78 = v65 == vc;
wire v79 = v78;
wire v7a = v25 & v79;
wire v91 = v7e == vc;
wire v92 = v91;
wire v93 = v28 & v92;
wire va7 = v61 | v7a | v93;
wire [31:0] vaa = ( va7 ) ? v4a : In_register_ESI;
wire [31:0] vc8 = vaa;
wire vca = vc8 == Out_register_ESI;
wire v112 = In_error_flag == Out_error_flag;
wire [31:0] v5 = 32'b00000000000000000000000000000101;
wire [31:0] v44 = ( v22 | v25 ) ? v5 : v5;
wire [31:0] v45 = In_register_EIP + v44;
wire [31:0] vd8 = v45;
wire vda = vd8 == Out_register_EIP;
wire v5c = v4c == vb;
wire v5d = v5c;
wire v5e = v22 & v5d;
wire v75 = v65 == vb;
wire v76 = v75;
wire v77 = v25 & v76;
wire v8e = v7e == vb;
wire v8f = v8e;
wire v90 = v28 & v8f;
wire va3 = v5e | v77 | v90;
wire [31:0] va6 = ( va3 ) ? v4a : In_register_EDX;
wire [31:0] vc4 = va6;
wire vc6 = vc4 == Out_register_EDX;
wire v62 = v4c == vd;
wire v63 = v62;
wire v64 = v22 & v63;
wire v7b = v65 == vd;
wire v7c = v7b;
wire v7d = v25 & v7c;
wire v94 = v7e == vd;
wire v95 = v94;
wire v96 = v28 & v95;
wire vaf = v64 | v7d | v96;
wire [31:0] vb2 = ( vaf ) ? v4a : In_register_ESP;
wire [31:0] vd0 = vb2;
wire vd2 = vd0 == Out_register_ESP;
wire [31:0] vdc = In_register_CSBASE;
wire vde = vdc == Out_register_CSBASE;
wire [31:0] ve0 = In_register_SSBASE;
wire ve2 = ve0 == Out_register_SSBASE;
wire [31:0] vec = In_register_GSBASE;
wire vee = vec == Out_register_GSBASE;
wire v59 = v4c == va;
wire v5a = v59;
wire v5b = v22 & v5a;
wire v72 = v65 == va;
wire v73 = v72;
wire v74 = v25 & v73;
wire v8b = v7e == va;
wire v8c = v8b;
wire v8d = v28 & v8c;
wire vab = v5b | v74 | v8d;
wire [31:0] vae = ( vab ) ? v4a : In_register_EDI;
wire [31:0] vcc = vae;
wire vce = vcc == Out_register_EDI;
wire [31:0] ve4 = In_register_ESBASE;
wire ve6 = ve4 == Out_register_ESBASE;
wire v105 = In_register_PF;
wire v107 = v105 == Out_register_PF;
wire [31:0] ve8 = In_register_DSBASE;
wire vea = ve8 == Out_register_DSBASE;
wire [7:0] vfc = In_register_DF;
wire vfe = vfc == Out_register_DF;
wire vff = vfe;
wire v4d = v4c == v6;
wire v4e = v4d;
wire v4f = v22 & v4e;
wire v66 = v65 == v6;
wire v67 = v66;
wire v68 = v25 & v67;
wire v7f = v7e == v6;
wire v80 = v7f;
wire v81 = v28 & v80;
wire v97 = v4f | v68 | v81;
wire [31:0] v9a = ( v97 ) ? v4a : In_register_EAX;
wire [31:0] vb8 = v9a;
wire vba = vb8 == Out_register_EAX;
wire [31:0] vf0 = In_register_FSBASE;
wire vf2 = vf0 == Out_register_FSBASE;
wire vf4 = In_register_AF;
wire vf6 = vf4 == Out_register_AF;
wire vf8 = In_register_CF;
wire vfa = vf8 == Out_register_CF;
wire v50 = v4c == v7;
wire v51 = v50;
wire v52 = v22 & v51;
wire v69 = v65 == v7;
wire v6a = v69;
wire v6b = v25 & v6a;
wire v82 = v7e == v7;
wire v83 = v82;
wire v84 = v28 & v83;
wire vb3 = v52 | v6b | v84;
wire [31:0] vb6 = ( vb3 ) ? v4a : In_register_EBP;
wire [31:0] vd4 = vb6;
wire vd6 = vd4 == Out_register_EBP;
wire v10d = In_register_ZF;
wire v10f = v10d == Out_register_ZF;
wire v113 = v2a & v103 & vbe & v10b & v1d & vc2 & vca & v112 & vda & vc6 & vd2 & vde & ve2 & vee & vce & ve6 & v107 & vea & vff & vba & vf2 & vf6 & vfa & vd6 & v10f;
wire v23b = v1ec | v23a | v113;
assign result = v23b;
endmodule
